-- ****************************************** --
-- * Integrated Systems Architecture        * --
-- * Lab 03: RISC-V                         * --  
-- * PACKAGE for TESTBENCH top-level RISC-V * --   
-- * Authors:                               * --
-- *  FIORAVANTI Simone S292612             * --
-- *  MOLINA Ottavio    S292527             * --
-- *  OTTINO Lorenzo    S281571             * --
-- ****************************************** --

package package_tb_RISC_V is
	constant PERIOD : time := 1 us;
	constant Nbit : positive := 32;
end package package_tb_RISC_V;
