package package_tb_RISC_V is
	constant PERIOD : time := 1 us;
	constant Nbit : positive := 32;
end package package_tb_RISC_V;
